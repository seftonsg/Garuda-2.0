module SCF_tb();
wire [63:0] o;
reg [63:0] i;
SCF SCF1(i, o);
integer i;
initial begin
 i= 16;

#10 
  $display ("Value of o is %d ",o);
end
endmodule
module SCF(i, o);
output [63:0] o;
reg [63:0] o;
input [63:0] i;
reg [63:0] internal0;
reg [63:0] internal1;
always @(*)
begin
 internal1 = 0;
 internal0 = 0;
 o = 0;
if ((((((((((i >> 26) & (-1 >> 58)) == 4) | ((((i >> 26) & (-1 >> 58)) == 1) & (((i >> 11) & (-1 >> 59)) == 1))) | ((((i >> 26) & (-1 >> 58)) == 7) & (((i >> 11) & (-1 >> 59)) == 0))) | ((((i >> 26) & (-1 >> 58)) == 6) & (((i >> 11) & (-1 >> 59)) == 0))) | ((((i >> 26) & (-1 >> 58)) == 1) & (((i >> 11) & (-1 >> 59)) == 0))) | (((i >> 26) & (-1 >> 58)) == 5)) | ((((((i >> 26) & (-1 >> 58)) == 0) & (((i >> 0) & (-1 >> 58)) == 9)) | ((((i >> 26) & (-1 >> 58)) == 0) & (((i >> 0) & (-1 >> 58)) == 8))) | ((((i >> 26) & (-1 >> 58)) == 2) | (((i >> 26) & (-1 >> 58)) == 3)))))
begin
if (~(((i >> 42) & (-1 >> 32)) == 0))
begin
 internal0 = i;
end
else begin
end
end
else begin
end
if (~(((((((((i >> 26) & (-1 >> 58)) == 4) | ((((i >> 26) & (-1 >> 58)) == 1) & (((i >> 11) & (-1 >> 59)) == 1))) | ((((i >> 26) & (-1 >> 58)) == 7) & (((i >> 11) & (-1 >> 59)) == 0))) | ((((i >> 26) & (-1 >> 58)) == 6) & (((i >> 11) & (-1 >> 59)) == 0))) | ((((i >> 26) & (-1 >> 58)) == 1) & (((i >> 11) & (-1 >> 59)) == 0))) | (((i >> 26) & (-1 >> 58)) == 5)) | ((((((i >> 26) & (-1 >> 58)) == 0) & (((i >> 0) & (-1 >> 58)) == 9)) | ((((i >> 26) & (-1 >> 58)) == 0) & (((i >> 0) & (-1 >> 58)) == 8))) | ((((i >> 26) & (-1 >> 58)) == 2) | (((i >> 26) & (-1 >> 58)) == 3)))))
begin
 internal1 = i;
end
else begin
end
 o = (internal0 | internal1);



end
endmodule

